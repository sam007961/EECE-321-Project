-- P321 Instruction Memory
-- Copyright (c) 2017 Mazen A. R. Saghir
-- Department of Electrical and Computer Engineering
-- American University of Beirut

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rom1024x32 is
  port (addr : in std_logic_vector(31 downto 0);
	data : out std_logic_vector(31 downto 0));
end entity;

architecture instrMem of rom1024x32 is
  type rom_array is array (0 to 45) of std_logic_vector (31 downto 0);
  constant rom: rom_array := (
"00111110100000000000000010010011",
"11111111110100000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"00000000010100000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"00000000110000000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"11111111110100000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"00000001001000000000000100010011",
"00000000001000001010000000100011",
"01000000100000000000000010010011",
"00000000010000000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"11111110100000000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"00000000011000000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"11111111011000000000000100010011",
"00000000001000001010000000100011",
"00000000010000001000000010010011",
"00000001100100000000000100010011",
"00000000001000001010000000100011",
"00111110100000000000000010010011",
"01000000100000000000000100010011",
"00000000000000000000001100110011",
"00000000000000000000001110110011",
"00000000010100111010010000010011",
"00000000000001000000100101100011",
"00000000000000001010000110000011",
"00000000000000010010001000000011",
"00000010010000011000001010110011", 
"00000000010100110000001100110011", 
"00000000010000001000000010010011",
"00000000010000010000000100010011",
"00000000000100111000001110010011",
"11111111111111101110000001101111", --corrected to -18
"00000000001100110001001100010011",
"00000000000000110000000001100111");
begin
  data <= rom(conv_integer(unsigned(addr(31 downto 2)))) when conv_integer(unsigned(addr(31 downto 0))) < 184 else "00000000000000000000000000000000";
end architecture;

